module sccb_timing_gen #(

) (
    
);

endmodule