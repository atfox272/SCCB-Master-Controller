module sccb_fsm #(

) (

);

endmodule